library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity Decoder_reg is
port (
i : in std_logic_vector ( 4 downto 0);
o : out std_logic_vector ( 31 downto 0)
);	
end Decoder_reg;

architecture Behavioral of Decoder_reg is
	SIGNAL sel: STD_LOGIC_VECTOR (31 DOWNTO 0) := (others => '0');




BEGIN
process (i)
BEGIN

o <= "11111111111111111111111111111111";
	if (i="00000") then o <= "00000000000000000000000000000001";
elsif (i="00001") then o <= "00000000000000000000000000000010";
elsif (i="00010") then o <= "00000000000000000000000000000100";
elsif (i="00011") then o <= "00000000000000000000000000001000";
elsif (i="00100") then o <= "00000000000000000000000000010000";
elsif (i="00101") then o <= "00000000000000000000000000100000";
elsif (i="00110") then o <= "00000000000000000000000001000000";
elsif (i="00111") then o <= "00000000000000000000000010000000";
elsif (i="01000") then o <= "00000000000000000000000100000000";
elsif (i="01001") then o <= "00000000000000000000001000000000";
elsif (i="01010") then o <= "00000000000000000000010000000000";
elsif (i="01011") then o <= "00000000000000000000100000000000";
elsif (i="01100") then o <= "00000000000000000001000000000000";
elsif (i="01101") then o <= "00000000000000000010000000000000";
elsif (i="01110") then o <= "00000000000000000100000000000000";
elsif (i="01111") then o <= "00000000000000001000000000000000";
elsif (i="10000") then o <= "00000000000000010000000000000000";
elsif (i="10001") then o <= "00000000000000100000000000000000";
elsif (i="10010") then o <= "00000000000001000000000000000000";
elsif (i="10011") then o <= "00000000000010000000000000000000";
elsif (i="10100") then o <= "00000000000100000000000000000000";
elsif (i="10101") then o <= "00000000001000000000000000000000";
elsif (i="10110") then o <= "00000000010000000000000000000000";
elsif (i="10111") then o <= "00000000100000000000000000000000";
elsif (i="11000") then o <= "00000001000000000000000000000000";
elsif (i="11001") then o <= "00000010000000000000000000000000";
elsif (i="11010") then o <= "00000100000000000000000000000000";
elsif (i="11011") then o <= "00001000000000000000000000000000";
elsif (i="11100") then o <= "00010000000000000000000000000000";
elsif (i="11101") then o <= "00100000000000000000000000000000";
elsif (i="11110") then o <= "01000000000000000000000000000000";
elsif (i="11111") then o <= "10000000000000000000000000000000";


end if;


end process;

end Behavioral;
